// layer_controller.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module layer_controller (
		input  wire        clk_clk,          //        clk.clk
		output wire [7:0]  leds_export,      //       leds.export
		output wire [8:0]  n1i1_export,      //       n1i1.export
		output wire [8:0]  n1i2_export,      //       n1i2.export
		output wire [8:0]  n1i3_export,      //       n1i3.export
		output wire [2:0]  n1ninputs_export, //  n1ninputs.export
		input  wire [8:0]  n1output_export,  //   n1output.export
		input  wire        n1ready_export,   //    n1ready.export
		output wire        n1start_export,   //    n1start.export
		output wire [16:0] n1w1_export,      //       n1w1.export
		output wire [16:0] n1w2_export,      //       n1w2.export
		output wire [16:0] n1w3_export,      //       n1w3.export
		input  wire        reset_reset,      //      reset.reset
		output wire        sdram_clk_clk,    //  sdram_clk.clk
		output wire [12:0] sdram_wire_addr,  // sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,    //           .ba
		output wire        sdram_wire_cas_n, //           .cas_n
		output wire        sdram_wire_cke,   //           .cke
		output wire        sdram_wire_cs_n,  //           .cs_n
		inout  wire [15:0] sdram_wire_dq,    //           .dq
		output wire [1:0]  sdram_wire_dqm,   //           .dqm
		output wire        sdram_wire_ras_n, //           .ras_n
		output wire        sdram_wire_we_n   //           .we_n
	);

	wire         clocks_sys_clk_clk;                                        // clocks:sys_clk_clk -> [cpu:clk, input_1_neuron_1:clk, input_2_neuron_1:clk, input_3_neuron_1:clk, irq_mapper:clk, jtag_uart:clk, leds:clk, mm_interconnect_0:clocks_sys_clk_clk, nInputs_neuron_1:clk, onchip_memory2_0:clk, output_neuron_1:clk, ready_neuron_1:clk, rst_controller:clk, sdram:clk, start_neuron_1:clk, weight_1_neuron_1:clk, weight_2_neuron_1:clk, weight_3_neuron_1:clk]
	wire  [31:0] cpu_data_master_readdata;                                  // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                               // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                               // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [26:0] cpu_data_master_address;                                   // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                      // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_write;                                     // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                 // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                           // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [26:0] cpu_instruction_master_address;                            // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                               // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;            // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;         // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;         // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;             // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;          // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;               // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;           // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;          // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;            // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [12:0] mm_interconnect_0_onchip_memory2_0_s1_address;             // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;          // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;               // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;           // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;               // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_leds_s1_chipselect;                      // mm_interconnect_0:leds_s1_chipselect -> leds:chipselect
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                        // leds:readdata -> mm_interconnect_0:leds_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                         // mm_interconnect_0:leds_s1_address -> leds:address
	wire         mm_interconnect_0_leds_s1_write;                           // mm_interconnect_0:leds_s1_write -> leds:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                       // mm_interconnect_0:leds_s1_writedata -> leds:writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                     // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                       // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                    // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [23:0] mm_interconnect_0_sdram_s1_address;                        // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                           // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                     // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                  // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                          // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                      // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_start_neuron_1_s1_chipselect;            // mm_interconnect_0:start_neuron_1_s1_chipselect -> start_neuron_1:chipselect
	wire  [31:0] mm_interconnect_0_start_neuron_1_s1_readdata;              // start_neuron_1:readdata -> mm_interconnect_0:start_neuron_1_s1_readdata
	wire   [1:0] mm_interconnect_0_start_neuron_1_s1_address;               // mm_interconnect_0:start_neuron_1_s1_address -> start_neuron_1:address
	wire         mm_interconnect_0_start_neuron_1_s1_write;                 // mm_interconnect_0:start_neuron_1_s1_write -> start_neuron_1:write_n
	wire  [31:0] mm_interconnect_0_start_neuron_1_s1_writedata;             // mm_interconnect_0:start_neuron_1_s1_writedata -> start_neuron_1:writedata
	wire         mm_interconnect_0_input_1_neuron_1_s1_chipselect;          // mm_interconnect_0:input_1_neuron_1_s1_chipselect -> input_1_neuron_1:chipselect
	wire  [31:0] mm_interconnect_0_input_1_neuron_1_s1_readdata;            // input_1_neuron_1:readdata -> mm_interconnect_0:input_1_neuron_1_s1_readdata
	wire   [1:0] mm_interconnect_0_input_1_neuron_1_s1_address;             // mm_interconnect_0:input_1_neuron_1_s1_address -> input_1_neuron_1:address
	wire         mm_interconnect_0_input_1_neuron_1_s1_write;               // mm_interconnect_0:input_1_neuron_1_s1_write -> input_1_neuron_1:write_n
	wire  [31:0] mm_interconnect_0_input_1_neuron_1_s1_writedata;           // mm_interconnect_0:input_1_neuron_1_s1_writedata -> input_1_neuron_1:writedata
	wire         mm_interconnect_0_input_2_neuron_1_s1_chipselect;          // mm_interconnect_0:input_2_neuron_1_s1_chipselect -> input_2_neuron_1:chipselect
	wire  [31:0] mm_interconnect_0_input_2_neuron_1_s1_readdata;            // input_2_neuron_1:readdata -> mm_interconnect_0:input_2_neuron_1_s1_readdata
	wire   [1:0] mm_interconnect_0_input_2_neuron_1_s1_address;             // mm_interconnect_0:input_2_neuron_1_s1_address -> input_2_neuron_1:address
	wire         mm_interconnect_0_input_2_neuron_1_s1_write;               // mm_interconnect_0:input_2_neuron_1_s1_write -> input_2_neuron_1:write_n
	wire  [31:0] mm_interconnect_0_input_2_neuron_1_s1_writedata;           // mm_interconnect_0:input_2_neuron_1_s1_writedata -> input_2_neuron_1:writedata
	wire         mm_interconnect_0_weight_1_neuron_1_s1_chipselect;         // mm_interconnect_0:weight_1_neuron_1_s1_chipselect -> weight_1_neuron_1:chipselect
	wire  [31:0] mm_interconnect_0_weight_1_neuron_1_s1_readdata;           // weight_1_neuron_1:readdata -> mm_interconnect_0:weight_1_neuron_1_s1_readdata
	wire   [1:0] mm_interconnect_0_weight_1_neuron_1_s1_address;            // mm_interconnect_0:weight_1_neuron_1_s1_address -> weight_1_neuron_1:address
	wire         mm_interconnect_0_weight_1_neuron_1_s1_write;              // mm_interconnect_0:weight_1_neuron_1_s1_write -> weight_1_neuron_1:write_n
	wire  [31:0] mm_interconnect_0_weight_1_neuron_1_s1_writedata;          // mm_interconnect_0:weight_1_neuron_1_s1_writedata -> weight_1_neuron_1:writedata
	wire         mm_interconnect_0_weight_2_neuron_1_s1_chipselect;         // mm_interconnect_0:weight_2_neuron_1_s1_chipselect -> weight_2_neuron_1:chipselect
	wire  [31:0] mm_interconnect_0_weight_2_neuron_1_s1_readdata;           // weight_2_neuron_1:readdata -> mm_interconnect_0:weight_2_neuron_1_s1_readdata
	wire   [1:0] mm_interconnect_0_weight_2_neuron_1_s1_address;            // mm_interconnect_0:weight_2_neuron_1_s1_address -> weight_2_neuron_1:address
	wire         mm_interconnect_0_weight_2_neuron_1_s1_write;              // mm_interconnect_0:weight_2_neuron_1_s1_write -> weight_2_neuron_1:write_n
	wire  [31:0] mm_interconnect_0_weight_2_neuron_1_s1_writedata;          // mm_interconnect_0:weight_2_neuron_1_s1_writedata -> weight_2_neuron_1:writedata
	wire  [31:0] mm_interconnect_0_output_neuron_1_s1_readdata;             // output_neuron_1:readdata -> mm_interconnect_0:output_neuron_1_s1_readdata
	wire   [1:0] mm_interconnect_0_output_neuron_1_s1_address;              // mm_interconnect_0:output_neuron_1_s1_address -> output_neuron_1:address
	wire  [31:0] mm_interconnect_0_ready_neuron_1_s1_readdata;              // ready_neuron_1:readdata -> mm_interconnect_0:ready_neuron_1_s1_readdata
	wire   [1:0] mm_interconnect_0_ready_neuron_1_s1_address;               // mm_interconnect_0:ready_neuron_1_s1_address -> ready_neuron_1:address
	wire         mm_interconnect_0_ninputs_neuron_1_s1_chipselect;          // mm_interconnect_0:nInputs_neuron_1_s1_chipselect -> nInputs_neuron_1:chipselect
	wire  [31:0] mm_interconnect_0_ninputs_neuron_1_s1_readdata;            // nInputs_neuron_1:readdata -> mm_interconnect_0:nInputs_neuron_1_s1_readdata
	wire   [1:0] mm_interconnect_0_ninputs_neuron_1_s1_address;             // mm_interconnect_0:nInputs_neuron_1_s1_address -> nInputs_neuron_1:address
	wire         mm_interconnect_0_ninputs_neuron_1_s1_write;               // mm_interconnect_0:nInputs_neuron_1_s1_write -> nInputs_neuron_1:write_n
	wire  [31:0] mm_interconnect_0_ninputs_neuron_1_s1_writedata;           // mm_interconnect_0:nInputs_neuron_1_s1_writedata -> nInputs_neuron_1:writedata
	wire         mm_interconnect_0_input_3_neuron_1_s1_chipselect;          // mm_interconnect_0:input_3_neuron_1_s1_chipselect -> input_3_neuron_1:chipselect
	wire  [31:0] mm_interconnect_0_input_3_neuron_1_s1_readdata;            // input_3_neuron_1:readdata -> mm_interconnect_0:input_3_neuron_1_s1_readdata
	wire   [1:0] mm_interconnect_0_input_3_neuron_1_s1_address;             // mm_interconnect_0:input_3_neuron_1_s1_address -> input_3_neuron_1:address
	wire         mm_interconnect_0_input_3_neuron_1_s1_write;               // mm_interconnect_0:input_3_neuron_1_s1_write -> input_3_neuron_1:write_n
	wire  [31:0] mm_interconnect_0_input_3_neuron_1_s1_writedata;           // mm_interconnect_0:input_3_neuron_1_s1_writedata -> input_3_neuron_1:writedata
	wire         mm_interconnect_0_weight_3_neuron_1_s1_chipselect;         // mm_interconnect_0:weight_3_neuron_1_s1_chipselect -> weight_3_neuron_1:chipselect
	wire  [31:0] mm_interconnect_0_weight_3_neuron_1_s1_readdata;           // weight_3_neuron_1:readdata -> mm_interconnect_0:weight_3_neuron_1_s1_readdata
	wire   [1:0] mm_interconnect_0_weight_3_neuron_1_s1_address;            // mm_interconnect_0:weight_3_neuron_1_s1_address -> weight_3_neuron_1:address
	wire         mm_interconnect_0_weight_3_neuron_1_s1_write;              // mm_interconnect_0:weight_3_neuron_1_s1_write -> weight_3_neuron_1:write_n
	wire  [31:0] mm_interconnect_0_weight_3_neuron_1_s1_writedata;          // mm_interconnect_0:weight_3_neuron_1_s1_writedata -> weight_3_neuron_1:writedata
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] cpu_irq_irq;                                               // irq_mapper:sender_irq -> cpu:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [cpu:reset_n, input_1_neuron_1:reset_n, input_2_neuron_1:reset_n, input_3_neuron_1:reset_n, irq_mapper:reset, jtag_uart:rst_n, leds:reset_n, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, nInputs_neuron_1:reset_n, onchip_memory2_0:reset, output_neuron_1:reset_n, ready_neuron_1:reset_n, rst_translator:in_reset, sdram:reset_n, start_neuron_1:reset_n, weight_1_neuron_1:reset_n, weight_2_neuron_1:reset_n, weight_3_neuron_1:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [cpu:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         cpu_debug_reset_request_reset;                             // cpu:debug_reset_request -> rst_controller:reset_in0
	wire         clocks_reset_source_reset;                                 // clocks:reset_source_reset -> rst_controller:reset_in1

	layer_controller_clocks clocks (
		.ref_clk_clk        (clk_clk),                   //      ref_clk.clk
		.ref_reset_reset    (reset_reset),               //    ref_reset.reset
		.sys_clk_clk        (clocks_sys_clk_clk),        //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),             //    sdram_clk.clk
		.reset_source_reset (clocks_reset_source_reset)  // reset_source.reset
	);

	layer_controller_cpu cpu (
		.clk                                 (clocks_sys_clk_clk),                                //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	layer_controller_input_1_neuron_1 input_1_neuron_1 (
		.clk        (clocks_sys_clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_input_1_neuron_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_input_1_neuron_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_input_1_neuron_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_input_1_neuron_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_input_1_neuron_1_s1_readdata),   //                    .readdata
		.out_port   (n1i1_export)                                       // external_connection.export
	);

	layer_controller_input_1_neuron_1 input_2_neuron_1 (
		.clk        (clocks_sys_clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_input_2_neuron_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_input_2_neuron_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_input_2_neuron_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_input_2_neuron_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_input_2_neuron_1_s1_readdata),   //                    .readdata
		.out_port   (n1i2_export)                                       // external_connection.export
	);

	layer_controller_input_1_neuron_1 input_3_neuron_1 (
		.clk        (clocks_sys_clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_input_3_neuron_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_input_3_neuron_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_input_3_neuron_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_input_3_neuron_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_input_3_neuron_1_s1_readdata),   //                    .readdata
		.out_port   (n1i3_export)                                       // external_connection.export
	);

	layer_controller_jtag_uart jtag_uart (
		.clk            (clocks_sys_clk_clk),                                        //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	layer_controller_leds leds (
		.clk        (clocks_sys_clk_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (leds_export)                           // external_connection.export
	);

	layer_controller_nInputs_neuron_1 ninputs_neuron_1 (
		.clk        (clocks_sys_clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_ninputs_neuron_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ninputs_neuron_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ninputs_neuron_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ninputs_neuron_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ninputs_neuron_1_s1_readdata),   //                    .readdata
		.out_port   (n1ninputs_export)                                  // external_connection.export
	);

	layer_controller_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clocks_sys_clk_clk),                               //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	layer_controller_output_neuron_1 output_neuron_1 (
		.clk      (clocks_sys_clk_clk),                            //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_0_output_neuron_1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_output_neuron_1_s1_readdata), //                    .readdata
		.in_port  (n1output_export)                                // external_connection.export
	);

	layer_controller_ready_neuron_1 ready_neuron_1 (
		.clk      (clocks_sys_clk_clk),                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address  (mm_interconnect_0_ready_neuron_1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_ready_neuron_1_s1_readdata), //                    .readdata
		.in_port  (n1ready_export)                                // external_connection.export
	);

	layer_controller_sdram sdram (
		.clk            (clocks_sys_clk_clk),                       //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	layer_controller_start_neuron_1 start_neuron_1 (
		.clk        (clocks_sys_clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_start_neuron_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_start_neuron_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_start_neuron_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_start_neuron_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_start_neuron_1_s1_readdata),   //                    .readdata
		.out_port   (n1start_export)                                  // external_connection.export
	);

	layer_controller_weight_1_neuron_1 weight_1_neuron_1 (
		.clk        (clocks_sys_clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (mm_interconnect_0_weight_1_neuron_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_weight_1_neuron_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_weight_1_neuron_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_weight_1_neuron_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_weight_1_neuron_1_s1_readdata),   //                    .readdata
		.out_port   (n1w1_export)                                        // external_connection.export
	);

	layer_controller_weight_1_neuron_1 weight_2_neuron_1 (
		.clk        (clocks_sys_clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (mm_interconnect_0_weight_2_neuron_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_weight_2_neuron_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_weight_2_neuron_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_weight_2_neuron_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_weight_2_neuron_1_s1_readdata),   //                    .readdata
		.out_port   (n1w2_export)                                        // external_connection.export
	);

	layer_controller_weight_1_neuron_1 weight_3_neuron_1 (
		.clk        (clocks_sys_clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (mm_interconnect_0_weight_3_neuron_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_weight_3_neuron_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_weight_3_neuron_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_weight_3_neuron_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_weight_3_neuron_1_s1_readdata),   //                    .readdata
		.out_port   (n1w3_export)                                        // external_connection.export
	);

	layer_controller_mm_interconnect_0 mm_interconnect_0 (
		.clocks_sys_clk_clk                      (clocks_sys_clk_clk),                                        //                  clocks_sys_clk.clk
		.cpu_reset_reset_bridge_in_reset_reset   (rst_controller_reset_out_reset),                            // cpu_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                 (cpu_data_master_address),                                   //                 cpu_data_master.address
		.cpu_data_master_waitrequest             (cpu_data_master_waitrequest),                               //                                .waitrequest
		.cpu_data_master_byteenable              (cpu_data_master_byteenable),                                //                                .byteenable
		.cpu_data_master_read                    (cpu_data_master_read),                                      //                                .read
		.cpu_data_master_readdata                (cpu_data_master_readdata),                                  //                                .readdata
		.cpu_data_master_write                   (cpu_data_master_write),                                     //                                .write
		.cpu_data_master_writedata               (cpu_data_master_writedata),                                 //                                .writedata
		.cpu_data_master_debugaccess             (cpu_data_master_debugaccess),                               //                                .debugaccess
		.cpu_instruction_master_address          (cpu_instruction_master_address),                            //          cpu_instruction_master.address
		.cpu_instruction_master_waitrequest      (cpu_instruction_master_waitrequest),                        //                                .waitrequest
		.cpu_instruction_master_read             (cpu_instruction_master_read),                               //                                .read
		.cpu_instruction_master_readdata         (cpu_instruction_master_readdata),                           //                                .readdata
		.cpu_debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),             //             cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),               //                                .write
		.cpu_debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),                //                                .read
		.cpu_debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),            //                                .readdata
		.cpu_debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),           //                                .writedata
		.cpu_debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),          //                                .byteenable
		.cpu_debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),         //                                .waitrequest
		.cpu_debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),         //                                .debugaccess
		.input_1_neuron_1_s1_address             (mm_interconnect_0_input_1_neuron_1_s1_address),             //             input_1_neuron_1_s1.address
		.input_1_neuron_1_s1_write               (mm_interconnect_0_input_1_neuron_1_s1_write),               //                                .write
		.input_1_neuron_1_s1_readdata            (mm_interconnect_0_input_1_neuron_1_s1_readdata),            //                                .readdata
		.input_1_neuron_1_s1_writedata           (mm_interconnect_0_input_1_neuron_1_s1_writedata),           //                                .writedata
		.input_1_neuron_1_s1_chipselect          (mm_interconnect_0_input_1_neuron_1_s1_chipselect),          //                                .chipselect
		.input_2_neuron_1_s1_address             (mm_interconnect_0_input_2_neuron_1_s1_address),             //             input_2_neuron_1_s1.address
		.input_2_neuron_1_s1_write               (mm_interconnect_0_input_2_neuron_1_s1_write),               //                                .write
		.input_2_neuron_1_s1_readdata            (mm_interconnect_0_input_2_neuron_1_s1_readdata),            //                                .readdata
		.input_2_neuron_1_s1_writedata           (mm_interconnect_0_input_2_neuron_1_s1_writedata),           //                                .writedata
		.input_2_neuron_1_s1_chipselect          (mm_interconnect_0_input_2_neuron_1_s1_chipselect),          //                                .chipselect
		.input_3_neuron_1_s1_address             (mm_interconnect_0_input_3_neuron_1_s1_address),             //             input_3_neuron_1_s1.address
		.input_3_neuron_1_s1_write               (mm_interconnect_0_input_3_neuron_1_s1_write),               //                                .write
		.input_3_neuron_1_s1_readdata            (mm_interconnect_0_input_3_neuron_1_s1_readdata),            //                                .readdata
		.input_3_neuron_1_s1_writedata           (mm_interconnect_0_input_3_neuron_1_s1_writedata),           //                                .writedata
		.input_3_neuron_1_s1_chipselect          (mm_interconnect_0_input_3_neuron_1_s1_chipselect),          //                                .chipselect
		.jtag_uart_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //     jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                .write
		.jtag_uart_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                .read
		.jtag_uart_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                .readdata
		.jtag_uart_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                .chipselect
		.leds_s1_address                         (mm_interconnect_0_leds_s1_address),                         //                         leds_s1.address
		.leds_s1_write                           (mm_interconnect_0_leds_s1_write),                           //                                .write
		.leds_s1_readdata                        (mm_interconnect_0_leds_s1_readdata),                        //                                .readdata
		.leds_s1_writedata                       (mm_interconnect_0_leds_s1_writedata),                       //                                .writedata
		.leds_s1_chipselect                      (mm_interconnect_0_leds_s1_chipselect),                      //                                .chipselect
		.nInputs_neuron_1_s1_address             (mm_interconnect_0_ninputs_neuron_1_s1_address),             //             nInputs_neuron_1_s1.address
		.nInputs_neuron_1_s1_write               (mm_interconnect_0_ninputs_neuron_1_s1_write),               //                                .write
		.nInputs_neuron_1_s1_readdata            (mm_interconnect_0_ninputs_neuron_1_s1_readdata),            //                                .readdata
		.nInputs_neuron_1_s1_writedata           (mm_interconnect_0_ninputs_neuron_1_s1_writedata),           //                                .writedata
		.nInputs_neuron_1_s1_chipselect          (mm_interconnect_0_ninputs_neuron_1_s1_chipselect),          //                                .chipselect
		.onchip_memory2_0_s1_address             (mm_interconnect_0_onchip_memory2_0_s1_address),             //             onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write               (mm_interconnect_0_onchip_memory2_0_s1_write),               //                                .write
		.onchip_memory2_0_s1_readdata            (mm_interconnect_0_onchip_memory2_0_s1_readdata),            //                                .readdata
		.onchip_memory2_0_s1_writedata           (mm_interconnect_0_onchip_memory2_0_s1_writedata),           //                                .writedata
		.onchip_memory2_0_s1_byteenable          (mm_interconnect_0_onchip_memory2_0_s1_byteenable),          //                                .byteenable
		.onchip_memory2_0_s1_chipselect          (mm_interconnect_0_onchip_memory2_0_s1_chipselect),          //                                .chipselect
		.onchip_memory2_0_s1_clken               (mm_interconnect_0_onchip_memory2_0_s1_clken),               //                                .clken
		.output_neuron_1_s1_address              (mm_interconnect_0_output_neuron_1_s1_address),              //              output_neuron_1_s1.address
		.output_neuron_1_s1_readdata             (mm_interconnect_0_output_neuron_1_s1_readdata),             //                                .readdata
		.ready_neuron_1_s1_address               (mm_interconnect_0_ready_neuron_1_s1_address),               //               ready_neuron_1_s1.address
		.ready_neuron_1_s1_readdata              (mm_interconnect_0_ready_neuron_1_s1_readdata),              //                                .readdata
		.sdram_s1_address                        (mm_interconnect_0_sdram_s1_address),                        //                        sdram_s1.address
		.sdram_s1_write                          (mm_interconnect_0_sdram_s1_write),                          //                                .write
		.sdram_s1_read                           (mm_interconnect_0_sdram_s1_read),                           //                                .read
		.sdram_s1_readdata                       (mm_interconnect_0_sdram_s1_readdata),                       //                                .readdata
		.sdram_s1_writedata                      (mm_interconnect_0_sdram_s1_writedata),                      //                                .writedata
		.sdram_s1_byteenable                     (mm_interconnect_0_sdram_s1_byteenable),                     //                                .byteenable
		.sdram_s1_readdatavalid                  (mm_interconnect_0_sdram_s1_readdatavalid),                  //                                .readdatavalid
		.sdram_s1_waitrequest                    (mm_interconnect_0_sdram_s1_waitrequest),                    //                                .waitrequest
		.sdram_s1_chipselect                     (mm_interconnect_0_sdram_s1_chipselect),                     //                                .chipselect
		.start_neuron_1_s1_address               (mm_interconnect_0_start_neuron_1_s1_address),               //               start_neuron_1_s1.address
		.start_neuron_1_s1_write                 (mm_interconnect_0_start_neuron_1_s1_write),                 //                                .write
		.start_neuron_1_s1_readdata              (mm_interconnect_0_start_neuron_1_s1_readdata),              //                                .readdata
		.start_neuron_1_s1_writedata             (mm_interconnect_0_start_neuron_1_s1_writedata),             //                                .writedata
		.start_neuron_1_s1_chipselect            (mm_interconnect_0_start_neuron_1_s1_chipselect),            //                                .chipselect
		.weight_1_neuron_1_s1_address            (mm_interconnect_0_weight_1_neuron_1_s1_address),            //            weight_1_neuron_1_s1.address
		.weight_1_neuron_1_s1_write              (mm_interconnect_0_weight_1_neuron_1_s1_write),              //                                .write
		.weight_1_neuron_1_s1_readdata           (mm_interconnect_0_weight_1_neuron_1_s1_readdata),           //                                .readdata
		.weight_1_neuron_1_s1_writedata          (mm_interconnect_0_weight_1_neuron_1_s1_writedata),          //                                .writedata
		.weight_1_neuron_1_s1_chipselect         (mm_interconnect_0_weight_1_neuron_1_s1_chipselect),         //                                .chipselect
		.weight_2_neuron_1_s1_address            (mm_interconnect_0_weight_2_neuron_1_s1_address),            //            weight_2_neuron_1_s1.address
		.weight_2_neuron_1_s1_write              (mm_interconnect_0_weight_2_neuron_1_s1_write),              //                                .write
		.weight_2_neuron_1_s1_readdata           (mm_interconnect_0_weight_2_neuron_1_s1_readdata),           //                                .readdata
		.weight_2_neuron_1_s1_writedata          (mm_interconnect_0_weight_2_neuron_1_s1_writedata),          //                                .writedata
		.weight_2_neuron_1_s1_chipselect         (mm_interconnect_0_weight_2_neuron_1_s1_chipselect),         //                                .chipselect
		.weight_3_neuron_1_s1_address            (mm_interconnect_0_weight_3_neuron_1_s1_address),            //            weight_3_neuron_1_s1.address
		.weight_3_neuron_1_s1_write              (mm_interconnect_0_weight_3_neuron_1_s1_write),              //                                .write
		.weight_3_neuron_1_s1_readdata           (mm_interconnect_0_weight_3_neuron_1_s1_readdata),           //                                .readdata
		.weight_3_neuron_1_s1_writedata          (mm_interconnect_0_weight_3_neuron_1_s1_writedata),          //                                .writedata
		.weight_3_neuron_1_s1_chipselect         (mm_interconnect_0_weight_3_neuron_1_s1_chipselect)          //                                .chipselect
	);

	layer_controller_irq_mapper irq_mapper (
		.clk           (clocks_sys_clk_clk),             //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (cpu_debug_reset_request_reset),      // reset_in0.reset
		.reset_in1      (clocks_reset_source_reset),          // reset_in1.reset
		.clk            (clocks_sys_clk_clk),                 //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
