library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity transfer_function is
	port(
		clk	: in std_logic;
		rst_n	: in std_logic;
		load	: in std_logic;
		input	: in std_logic_vector(16 downto 0);
		y		: out std_logic_vector(8 downto 0);
		eop	: out std_logic									-- end of process
	);
end entity transfer_function;

architecture transfer_function_behaviour of transfer_function is
	signal x : std_logic_vector(10 downto 0);
begin
	transfer: process(clk, rst_n) is
	begin
		if rst_n = '0' then
			x <= (others => '0');
		elsif rising_edge(clk)then
		--else
			if signed(input) <= -768 then								-- 11111110100000000	 in fixed point is this -3
				y <= "100000000";
			elsif signed(input) >= 768 then							-- 00000001100000000	 in fixed point is this 3
				y <= "011111111";
			else
				x <= input(16) & input(9 downto 0);
				case x is 
					when "10100000000" => y <= "100000010";
					when "10100000001" => y <= "100000010";
					when "10100000010" => y <= "100000010";
					when "10100000011" => y <= "100000010";
					when "10100000100" => y <= "100000010";
					when "10100000101" => y <= "100000010";
					when "10100000110" => y <= "100000010";
					when "10100000111" => y <= "100000010";
					when "10100001000" => y <= "100000010";
					when "10100001001" => y <= "100000010";
					when "10100001010" => y <= "100000010";
					when "10100001011" => y <= "100000010";
					when "10100001100" => y <= "100000010";
					when "10100001101" => y <= "100000010";
					when "10100001110" => y <= "100000010";
					when "10100001111" => y <= "100000010";
					when "10100010000" => y <= "100000010";
					when "10100010001" => y <= "100000010";
					when "10100010010" => y <= "100000010";
					when "10100010011" => y <= "100000010";
					when "10100010100" => y <= "100000010";
					when "10100010101" => y <= "100000010";
					when "10100010110" => y <= "100000010";
					when "10100010111" => y <= "100000010";
					when "10100011000" => y <= "100000010";
					when "10100011001" => y <= "100000010";
					when "10100011010" => y <= "100000010";
					when "10100011011" => y <= "100000010";
					when "10100011100" => y <= "100000010";
					when "10100011101" => y <= "100000010";
					when "10100011110" => y <= "100000010";
					when "10100011111" => y <= "100000010";
					when "10100100000" => y <= "100000010";
					when "10100100001" => y <= "100000010";
					when "10100100010" => y <= "100000010";
					when "10100100011" => y <= "100000010";
					when "10100100100" => y <= "100000010";
					when "10100100101" => y <= "100000010";
					when "10100100110" => y <= "100000010";
					when "10100100111" => y <= "100000010";
					when "10100101000" => y <= "100000010";
					when "10100101001" => y <= "100000010";
					when "10100101010" => y <= "100000010";
					when "10100101011" => y <= "100000010";
					when "10100101100" => y <= "100000010";
					when "10100101101" => y <= "100000010";
					when "10100101110" => y <= "100000010";
					when "10100101111" => y <= "100000010";
					when "10100110000" => y <= "100000010";
					when "10100110001" => y <= "100000010";
					when "10100110010" => y <= "100000010";
					when "10100110011" => y <= "100000010";
					when "10100110100" => y <= "100000010";
					when "10100110101" => y <= "100000010";
					when "10100110110" => y <= "100000010";
					when "10100110111" => y <= "100000010";
					when "10100111000" => y <= "100000010";
					when "10100111001" => y <= "100000010";
					when "10100111010" => y <= "100000010";
					when "10100111011" => y <= "100000011";
					when "10100111100" => y <= "100000011";
					when "10100111101" => y <= "100000011";
					when "10100111110" => y <= "100000011";
					when "10100111111" => y <= "100000011";
					when "10101000000" => y <= "100000011";
					when "10101000001" => y <= "100000011";
					when "10101000010" => y <= "100000011";
					when "10101000011" => y <= "100000011";
					when "10101000100" => y <= "100000011";
					when "10101000101" => y <= "100000011";
					when "10101000110" => y <= "100000011";
					when "10101000111" => y <= "100000011";
					when "10101001000" => y <= "100000011";
					when "10101001001" => y <= "100000011";
					when "10101001010" => y <= "100000011";
					when "10101001011" => y <= "100000011";
					when "10101001100" => y <= "100000011";
					when "10101001101" => y <= "100000011";
					when "10101001110" => y <= "100000011";
					when "10101001111" => y <= "100000011";
					when "10101010000" => y <= "100000011";
					when "10101010001" => y <= "100000011";
					when "10101010010" => y <= "100000011";
					when "10101010011" => y <= "100000011";
					when "10101010100" => y <= "100000011";
					when "10101010101" => y <= "100000011";
					when "10101010110" => y <= "100000011";
					when "10101010111" => y <= "100000011";
					when "10101011000" => y <= "100000011";
					when "10101011001" => y <= "100000011";
					when "10101011010" => y <= "100000011";
					when "10101011011" => y <= "100000011";
					when "10101011100" => y <= "100000011";
					when "10101011101" => y <= "100000011";
					when "10101011110" => y <= "100000011";
					when "10101011111" => y <= "100000011";
					when "10101100000" => y <= "100000011";
					when "10101100001" => y <= "100000011";
					when "10101100010" => y <= "100000011";
					when "10101100011" => y <= "100000011";
					when "10101100100" => y <= "100000011";
					when "10101100101" => y <= "100000011";
					when "10101100110" => y <= "100000011";
					when "10101100111" => y <= "100000011";
					when "10101101000" => y <= "100000011";
					when "10101101001" => y <= "100000011";
					when "10101101010" => y <= "100000011";
					when "10101101011" => y <= "100000011";
					when "10101101100" => y <= "100000011";
					when "10101101101" => y <= "100000011";
					when "10101101110" => y <= "100000011";
					when "10101101111" => y <= "100000100";
					when "10101110000" => y <= "100000100";
					when "10101110001" => y <= "100000100";
					when "10101110010" => y <= "100000100";
					when "10101110011" => y <= "100000100";
					when "10101110100" => y <= "100000100";
					when "10101110101" => y <= "100000100";
					when "10101110110" => y <= "100000100";
					when "10101110111" => y <= "100000100";
					when "10101111000" => y <= "100000100";
					when "10101111001" => y <= "100000100";
					when "10101111010" => y <= "100000100";
					when "10101111011" => y <= "100000100";
					when "10101111100" => y <= "100000100";
					when "10101111101" => y <= "100000100";
					when "10101111110" => y <= "100000100";
					when "10101111111" => y <= "100000100";
					when "10110000000" => y <= "100000100";
					when "10110000001" => y <= "100000100";
					when "10110000010" => y <= "100000100";
					when "10110000011" => y <= "100000100";
					when "10110000100" => y <= "100000100";
					when "10110000101" => y <= "100000100";
					when "10110000110" => y <= "100000100";
					when "10110000111" => y <= "100000100";
					when "10110001000" => y <= "100000100";
					when "10110001001" => y <= "100000100";
					when "10110001010" => y <= "100000100";
					when "10110001011" => y <= "100000100";
					when "10110001100" => y <= "100000100";
					when "10110001101" => y <= "100000100";
					when "10110001110" => y <= "100000100";
					when "10110001111" => y <= "100000100";
					when "10110010000" => y <= "100000100";
					when "10110010001" => y <= "100000100";
					when "10110010010" => y <= "100000100";
					when "10110010011" => y <= "100000100";
					when "10110010100" => y <= "100000101";
					when "10110010101" => y <= "100000101";
					when "10110010110" => y <= "100000101";
					when "10110010111" => y <= "100000101";
					when "10110011000" => y <= "100000101";
					when "10110011001" => y <= "100000101";
					when "10110011010" => y <= "100000101";
					when "10110011011" => y <= "100000101";
					when "10110011100" => y <= "100000101";
					when "10110011101" => y <= "100000101";
					when "10110011110" => y <= "100000101";
					when "10110011111" => y <= "100000101";
					when "10110100000" => y <= "100000101";
					when "10110100001" => y <= "100000101";
					when "10110100010" => y <= "100000101";
					when "10110100011" => y <= "100000101";
					when "10110100100" => y <= "100000101";
					when "10110100101" => y <= "100000101";
					when "10110100110" => y <= "100000101";
					when "10110100111" => y <= "100000101";
					when "10110101000" => y <= "100000101";
					when "10110101001" => y <= "100000101";
					when "10110101010" => y <= "100000101";
					when "10110101011" => y <= "100000101";
					when "10110101100" => y <= "100000101";
					when "10110101101" => y <= "100000101";
					when "10110101110" => y <= "100000101";
					when "10110101111" => y <= "100000101";
					when "10110110000" => y <= "100000101";
					when "10110110001" => y <= "100000110";
					when "10110110010" => y <= "100000110";
					when "10110110011" => y <= "100000110";
					when "10110110100" => y <= "100000110";
					when "10110110101" => y <= "100000110";
					when "10110110110" => y <= "100000110";
					when "10110110111" => y <= "100000110";
					when "10110111000" => y <= "100000110";
					when "10110111001" => y <= "100000110";
					when "10110111010" => y <= "100000110";
					when "10110111011" => y <= "100000110";
					when "10110111100" => y <= "100000110";
					when "10110111101" => y <= "100000110";
					when "10110111110" => y <= "100000110";
					when "10110111111" => y <= "100000110";
					when "10111000000" => y <= "100000110";
					when "10111000001" => y <= "100000110";
					when "10111000010" => y <= "100000110";
					when "10111000011" => y <= "100000110";
					when "10111000100" => y <= "100000110";
					when "10111000101" => y <= "100000110";
					when "10111000110" => y <= "100000110";
					when "10111000111" => y <= "100000110";
					when "10111001000" => y <= "100000110";
					when "10111001001" => y <= "100000111";
					when "10111001010" => y <= "100000111";
					when "10111001011" => y <= "100000111";
					when "10111001100" => y <= "100000111";
					when "10111001101" => y <= "100000111";
					when "10111001110" => y <= "100000111";
					when "10111001111" => y <= "100000111";
					when "10111010000" => y <= "100000111";
					when "10111010001" => y <= "100000111";
					when "10111010010" => y <= "100000111";
					when "10111010011" => y <= "100000111";
					when "10111010100" => y <= "100000111";
					when "10111010101" => y <= "100000111";
					when "10111010110" => y <= "100000111";
					when "10111010111" => y <= "100000111";
					when "10111011000" => y <= "100000111";
					when "10111011001" => y <= "100000111";
					when "10111011010" => y <= "100000111";
					when "10111011011" => y <= "100000111";
					when "10111011100" => y <= "100000111";
					when "10111011101" => y <= "100001000";
					when "10111011110" => y <= "100001000";
					when "10111011111" => y <= "100001000";
					when "10111100000" => y <= "100001000";
					when "10111100001" => y <= "100001000";
					when "10111100010" => y <= "100001000";
					when "10111100011" => y <= "100001000";
					when "10111100100" => y <= "100001000";
					when "10111100101" => y <= "100001000";
					when "10111100110" => y <= "100001000";
					when "10111100111" => y <= "100001000";
					when "10111101000" => y <= "100001000";
					when "10111101001" => y <= "100001000";
					when "10111101010" => y <= "100001000";
					when "10111101011" => y <= "100001000";
					when "10111101100" => y <= "100001000";
					when "10111101101" => y <= "100001000";
					when "10111101110" => y <= "100001001";
					when "10111101111" => y <= "100001001";
					when "10111110000" => y <= "100001001";
					when "10111110001" => y <= "100001001";
					when "10111110010" => y <= "100001001";
					when "10111110011" => y <= "100001001";
					when "10111110100" => y <= "100001001";
					when "10111110101" => y <= "100001001";
					when "10111110110" => y <= "100001001";
					when "10111110111" => y <= "100001001";
					when "10111111000" => y <= "100001001";
					when "10111111001" => y <= "100001001";
					when "10111111010" => y <= "100001001";
					when "10111111011" => y <= "100001001";
					when "10111111100" => y <= "100001001";
					when "10111111101" => y <= "100001001";
					when "10111111110" => y <= "100001010";
					when "10111111111" => y <= "100001010";
					when "11000000000" => y <= "100001010";
					when "11000000001" => y <= "100001010";
					when "11000000010" => y <= "100001010";
					when "11000000011" => y <= "100001010";
					when "11000000100" => y <= "100001010";
					when "11000000101" => y <= "100001010";
					when "11000000110" => y <= "100001010";
					when "11000000111" => y <= "100001010";
					when "11000001000" => y <= "100001010";
					when "11000001001" => y <= "100001010";
					when "11000001010" => y <= "100001010";
					when "11000001011" => y <= "100001011";
					when "11000001100" => y <= "100001011";
					when "11000001101" => y <= "100001011";
					when "11000001110" => y <= "100001011";
					when "11000001111" => y <= "100001011";
					when "11000010000" => y <= "100001011";
					when "11000010001" => y <= "100001011";
					when "11000010010" => y <= "100001011";
					when "11000010011" => y <= "100001011";
					when "11000010100" => y <= "100001011";
					when "11000010101" => y <= "100001011";
					when "11000010110" => y <= "100001011";
					when "11000010111" => y <= "100001011";
					when "11000011000" => y <= "100001100";
					when "11000011001" => y <= "100001100";
					when "11000011010" => y <= "100001100";
					when "11000011011" => y <= "100001100";
					when "11000011100" => y <= "100001100";
					when "11000011101" => y <= "100001100";
					when "11000011110" => y <= "100001100";
					when "11000011111" => y <= "100001100";
					when "11000100000" => y <= "100001100";
					when "11000100001" => y <= "100001100";
					when "11000100010" => y <= "100001100";
					when "11000100011" => y <= "100001101";
					when "11000100100" => y <= "100001101";
					when "11000100101" => y <= "100001101";
					when "11000100110" => y <= "100001101";
					when "11000100111" => y <= "100001101";
					when "11000101000" => y <= "100001101";
					when "11000101001" => y <= "100001101";
					when "11000101010" => y <= "100001101";
					when "11000101011" => y <= "100001101";
					when "11000101100" => y <= "100001101";
					when "11000101101" => y <= "100001101";
					when "11000101110" => y <= "100001110";
					when "11000101111" => y <= "100001110";
					when "11000110000" => y <= "100001110";
					when "11000110001" => y <= "100001110";
					when "11000110010" => y <= "100001110";
					when "11000110011" => y <= "100001110";
					when "11000110100" => y <= "100001110";
					when "11000110101" => y <= "100001110";
					when "11000110110" => y <= "100001110";
					when "11000110111" => y <= "100001111";
					when "11000111000" => y <= "100001111";
					when "11000111001" => y <= "100001111";
					when "11000111010" => y <= "100001111";
					when "11000111011" => y <= "100001111";
					when "11000111100" => y <= "100001111";
					when "11000111101" => y <= "100001111";
					when "11000111110" => y <= "100001111";
					when "11000111111" => y <= "100001111";
					when "11001000000" => y <= "100010000";
					when "11001000001" => y <= "100010000";
					when "11001000010" => y <= "100010000";
					when "11001000011" => y <= "100010000";
					when "11001000100" => y <= "100010000";
					when "11001000101" => y <= "100010000";
					when "11001000110" => y <= "100010000";
					when "11001000111" => y <= "100010000";
					when "11001001000" => y <= "100010000";
					when "11001001001" => y <= "100010001";
					when "11001001010" => y <= "100010001";
					when "11001001011" => y <= "100010001";
					when "11001001100" => y <= "100010001";
					when "11001001101" => y <= "100010001";
					when "11001001110" => y <= "100010001";
					when "11001001111" => y <= "100010001";
					when "11001010000" => y <= "100010001";
					when "11001010001" => y <= "100010010";
					when "11001010010" => y <= "100010010";
					when "11001010011" => y <= "100010010";
					when "11001010100" => y <= "100010010";
					when "11001010101" => y <= "100010010";
					when "11001010110" => y <= "100010010";
					when "11001010111" => y <= "100010010";
					when "11001011000" => y <= "100010010";
					when "11001011001" => y <= "100010011";
					when "11001011010" => y <= "100010011";
					when "11001011011" => y <= "100010011";
					when "11001011100" => y <= "100010011";
					when "11001011101" => y <= "100010011";
					when "11001011110" => y <= "100010011";
					when "11001011111" => y <= "100010011";
					when "11001100000" => y <= "100010100";
					when "11001100001" => y <= "100010100";
					when "11001100010" => y <= "100010100";
					when "11001100011" => y <= "100010100";
					when "11001100100" => y <= "100010100";
					when "11001100101" => y <= "100010100";
					when "11001100110" => y <= "100010100";
					when "11001100111" => y <= "100010101";
					when "11001101000" => y <= "100010101";
					when "11001101001" => y <= "100010101";
					when "11001101010" => y <= "100010101";
					when "11001101011" => y <= "100010101";
					when "11001101100" => y <= "100010101";
					when "11001101101" => y <= "100010110";
					when "11001101110" => y <= "100010110";
					when "11001101111" => y <= "100010110";
					when "11001110000" => y <= "100010110";
					when "11001110001" => y <= "100010110";
					when "11001110010" => y <= "100010110";
					when "11001110011" => y <= "100010111";
					when "11001110100" => y <= "100010111";
					when "11001110101" => y <= "100010111";
					when "11001110110" => y <= "100010111";
					when "11001110111" => y <= "100010111";
					when "11001111000" => y <= "100010111";
					when "11001111001" => y <= "100011000";
					when "11001111010" => y <= "100011000";
					when "11001111011" => y <= "100011000";
					when "11001111100" => y <= "100011000";
					when "11001111101" => y <= "100011000";
					when "11001111110" => y <= "100011000";
					when "11001111111" => y <= "100011001";
					when "11010000000" => y <= "100011001";
					when "11010000001" => y <= "100011001";
					when "11010000010" => y <= "100011001";
					when "11010000011" => y <= "100011001";
					when "11010000100" => y <= "100011010";
					when "11010000101" => y <= "100011010";
					when "11010000110" => y <= "100011010";
					when "11010000111" => y <= "100011010";
					when "11010001000" => y <= "100011010";
					when "11010001001" => y <= "100011010";
					when "11010001010" => y <= "100011011";
					when "11010001011" => y <= "100011011";
					when "11010001100" => y <= "100011011";
					when "11010001101" => y <= "100011011";
					when "11010001110" => y <= "100011011";
					when "11010001111" => y <= "100011100";
					when "11010010000" => y <= "100011100";
					when "11010010001" => y <= "100011100";
					when "11010010010" => y <= "100011100";
					when "11010010011" => y <= "100011100";
					when "11010010100" => y <= "100011101";
					when "11010010101" => y <= "100011101";
					when "11010010110" => y <= "100011101";
					when "11010010111" => y <= "100011101";
					when "11010011000" => y <= "100011110";
					when "11010011001" => y <= "100011110";
					when "11010011010" => y <= "100011110";
					when "11010011011" => y <= "100011110";
					when "11010011100" => y <= "100011110";
					when "11010011101" => y <= "100011111";
					when "11010011110" => y <= "100011111";
					when "11010011111" => y <= "100011111";
					when "11010100000" => y <= "100011111";
					when "11010100001" => y <= "100011111";
					when "11010100010" => y <= "100100000";
					when "11010100011" => y <= "100100000";
					when "11010100100" => y <= "100100000";
					when "11010100101" => y <= "100100000";
					when "11010100110" => y <= "100100001";
					when "11010100111" => y <= "100100001";
					when "11010101000" => y <= "100100001";
					when "11010101001" => y <= "100100001";
					when "11010101010" => y <= "100100010";
					when "11010101011" => y <= "100100010";
					when "11010101100" => y <= "100100010";
					when "11010101101" => y <= "100100010";
					when "11010101110" => y <= "100100011";
					when "11010101111" => y <= "100100011";
					when "11010110000" => y <= "100100011";
					when "11010110001" => y <= "100100011";
					when "11010110010" => y <= "100100100";
					when "11010110011" => y <= "100100100";
					when "11010110100" => y <= "100100100";
					when "11010110101" => y <= "100100100";
					when "11010110110" => y <= "100100101";
					when "11010110111" => y <= "100100101";
					when "11010111000" => y <= "100100101";
					when "11010111001" => y <= "100100101";
					when "11010111010" => y <= "100100110";
					when "11010111011" => y <= "100100110";
					when "11010111100" => y <= "100100110";
					when "11010111101" => y <= "100100111";
					when "11010111110" => y <= "100100111";
					when "11010111111" => y <= "100100111";
					when "11011000000" => y <= "100100111";
					when "11011000001" => y <= "100101000";
					when "11011000010" => y <= "100101000";
					when "11011000011" => y <= "100101000";
					when "11011000100" => y <= "100101000";
					when "11011000101" => y <= "100101001";
					when "11011000110" => y <= "100101001";
					when "11011000111" => y <= "100101001";
					when "11011001000" => y <= "100101010";
					when "11011001001" => y <= "100101010";
					when "11011001010" => y <= "100101010";
					when "11011001011" => y <= "100101011";
					when "11011001100" => y <= "100101011";
					when "11011001101" => y <= "100101011";
					when "11011001110" => y <= "100101011";
					when "11011001111" => y <= "100101100";
					when "11011010000" => y <= "100101100";
					when "11011010001" => y <= "100101100";
					when "11011010010" => y <= "100101101";
					when "11011010011" => y <= "100101101";
					when "11011010100" => y <= "100101101";
					when "11011010101" => y <= "100101110";
					when "11011010110" => y <= "100101110";
					when "11011010111" => y <= "100101110";
					when "11011011000" => y <= "100101111";
					when "11011011001" => y <= "100101111";
					when "11011011010" => y <= "100101111";
					when "11011011011" => y <= "100110000";
					when "11011011100" => y <= "100110000";
					when "11011011101" => y <= "100110000";
					when "11011011110" => y <= "100110001";
					when "11011011111" => y <= "100110001";
					when "11011100000" => y <= "100110001";
					when "11011100001" => y <= "100110010";
					when "11011100010" => y <= "100110010";
					when "11011100011" => y <= "100110010";
					when "11011100100" => y <= "100110011";
					when "11011100101" => y <= "100110011";
					when "11011100110" => y <= "100110011";
					when "11011100111" => y <= "100110100";
					when "11011101000" => y <= "100110100";
					when "11011101001" => y <= "100110101";
					when "11011101010" => y <= "100110101";
					when "11011101011" => y <= "100110101";
					when "11011101100" => y <= "100110110";
					when "11011101101" => y <= "100110110";
					when "11011101110" => y <= "100110110";
					when "11011101111" => y <= "100110111";
					when "11011110000" => y <= "100110111";
					when "11011110001" => y <= "100111000";
					when "11011110010" => y <= "100111000";
					when "11011110011" => y <= "100111000";
					when "11011110100" => y <= "100111001";
					when "11011110101" => y <= "100111001";
					when "11011110110" => y <= "100111001";
					when "11011110111" => y <= "100111010";
					when "11011111000" => y <= "100111010";
					when "11011111001" => y <= "100111011";
					when "11011111010" => y <= "100111011";
					when "11011111011" => y <= "100111011";
					when "11011111100" => y <= "100111100";
					when "11011111101" => y <= "100111100";
					when "11011111110" => y <= "100111101";
					when "11011111111" => y <= "100111101";
					when "11100000000" => y <= "100111110";
					when "11100000001" => y <= "100111110";
					when "11100000010" => y <= "100111110";
					when "11100000011" => y <= "100111111";
					when "11100000100" => y <= "100111111";
					when "11100000101" => y <= "101000000";
					when "11100000110" => y <= "101000000";
					when "11100000111" => y <= "101000001";
					when "11100001000" => y <= "101000001";
					when "11100001001" => y <= "101000001";
					when "11100001010" => y <= "101000010";
					when "11100001011" => y <= "101000010";
					when "11100001100" => y <= "101000011";
					when "11100001101" => y <= "101000011";
					when "11100001110" => y <= "101000100";
					when "11100001111" => y <= "101000100";
					when "11100010000" => y <= "101000101";
					when "11100010001" => y <= "101000101";
					when "11100010010" => y <= "101000110";
					when "11100010011" => y <= "101000110";
					when "11100010100" => y <= "101000110";
					when "11100010101" => y <= "101000111";
					when "11100010110" => y <= "101000111";
					when "11100010111" => y <= "101001000";
					when "11100011000" => y <= "101001000";
					when "11100011001" => y <= "101001001";
					when "11100011010" => y <= "101001001";
					when "11100011011" => y <= "101001010";
					when "11100011100" => y <= "101001010";
					when "11100011101" => y <= "101001011";
					when "11100011110" => y <= "101001011";
					when "11100011111" => y <= "101001100";
					when "11100100000" => y <= "101001100";
					when "11100100001" => y <= "101001101";
					when "11100100010" => y <= "101001101";
					when "11100100011" => y <= "101001110";
					when "11100100100" => y <= "101001110";
					when "11100100101" => y <= "101001111";
					when "11100100110" => y <= "101001111";
					when "11100100111" => y <= "101010000";
					when "11100101000" => y <= "101010000";
					when "11100101001" => y <= "101010001";
					when "11100101010" => y <= "101010001";
					when "11100101011" => y <= "101010010";
					when "11100101100" => y <= "101010011";
					when "11100101101" => y <= "101010011";
					when "11100101110" => y <= "101010100";
					when "11100101111" => y <= "101010100";
					when "11100110000" => y <= "101010101";
					when "11100110001" => y <= "101010101";
					when "11100110010" => y <= "101010110";
					when "11100110011" => y <= "101010110";
					when "11100110100" => y <= "101010111";
					when "11100110101" => y <= "101011000";
					when "11100110110" => y <= "101011000";
					when "11100110111" => y <= "101011001";
					when "11100111000" => y <= "101011001";
					when "11100111001" => y <= "101011010";
					when "11100111010" => y <= "101011010";
					when "11100111011" => y <= "101011011";
					when "11100111100" => y <= "101011100";
					when "11100111101" => y <= "101011100";
					when "11100111110" => y <= "101011101";
					when "11100111111" => y <= "101011101";
					when "11101000000" => y <= "101011110";
					when "11101000001" => y <= "101011110";
					when "11101000010" => y <= "101011111";
					when "11101000011" => y <= "101100000";
					when "11101000100" => y <= "101100000";
					when "11101000101" => y <= "101100001";
					when "11101000110" => y <= "101100010";
					when "11101000111" => y <= "101100010";
					when "11101001000" => y <= "101100011";
					when "11101001001" => y <= "101100011";
					when "11101001010" => y <= "101100100";
					when "11101001011" => y <= "101100101";
					when "11101001100" => y <= "101100101";
					when "11101001101" => y <= "101100110";
					when "11101001110" => y <= "101100111";
					when "11101001111" => y <= "101100111";
					when "11101010000" => y <= "101101000";
					when "11101010001" => y <= "101101000";
					when "11101010010" => y <= "101101001";
					when "11101010011" => y <= "101101010";
					when "11101010100" => y <= "101101010";
					when "11101010101" => y <= "101101011";
					when "11101010110" => y <= "101101100";
					when "11101010111" => y <= "101101100";
					when "11101011000" => y <= "101101101";
					when "11101011001" => y <= "101101110";
					when "11101011010" => y <= "101101110";
					when "11101011011" => y <= "101101111";
					when "11101011100" => y <= "101110000";
					when "11101011101" => y <= "101110000";
					when "11101011110" => y <= "101110001";
					when "11101011111" => y <= "101110010";
					when "11101100000" => y <= "101110011";
					when "11101100001" => y <= "101110011";
					when "11101100010" => y <= "101110100";
					when "11101100011" => y <= "101110101";
					when "11101100100" => y <= "101110101";
					when "11101100101" => y <= "101110110";
					when "11101100110" => y <= "101110111";
					when "11101100111" => y <= "101110111";
					when "11101101000" => y <= "101111000";
					when "11101101001" => y <= "101111001";
					when "11101101010" => y <= "101111010";
					when "11101101011" => y <= "101111010";
					when "11101101100" => y <= "101111011";
					when "11101101101" => y <= "101111100";
					when "11101101110" => y <= "101111101";
					when "11101101111" => y <= "101111101";
					when "11101110000" => y <= "101111110";
					when "11101110001" => y <= "101111111";
					when "11101110010" => y <= "101111111";
					when "11101110011" => y <= "110000000";
					when "11101110100" => y <= "110000001";
					when "11101110101" => y <= "110000010";
					when "11101110110" => y <= "110000010";
					when "11101110111" => y <= "110000011";
					when "11101111000" => y <= "110000100";
					when "11101111001" => y <= "110000101";
					when "11101111010" => y <= "110000110";
					when "11101111011" => y <= "110000110";
					when "11101111100" => y <= "110000111";
					when "11101111101" => y <= "110001000";
					when "11101111110" => y <= "110001001";
					when "11101111111" => y <= "110001001";
					when "11110000000" => y <= "110001010";
					when "11110000001" => y <= "110001011";
					when "11110000010" => y <= "110001100";
					when "11110000011" => y <= "110001101";
					when "11110000100" => y <= "110001101";
					when "11110000101" => y <= "110001110";
					when "11110000110" => y <= "110001111";
					when "11110000111" => y <= "110010000";
					when "11110001000" => y <= "110010001";
					when "11110001001" => y <= "110010001";
					when "11110001010" => y <= "110010010";
					when "11110001011" => y <= "110010011";
					when "11110001100" => y <= "110010100";
					when "11110001101" => y <= "110010101";
					when "11110001110" => y <= "110010101";
					when "11110001111" => y <= "110010110";
					when "11110010000" => y <= "110010111";
					when "11110010001" => y <= "110011000";
					when "11110010010" => y <= "110011001";
					when "11110010011" => y <= "110011010";
					when "11110010100" => y <= "110011010";
					when "11110010101" => y <= "110011011";
					when "11110010110" => y <= "110011100";
					when "11110010111" => y <= "110011101";
					when "11110011000" => y <= "110011110";
					when "11110011001" => y <= "110011111";
					when "11110011010" => y <= "110100000";
					when "11110011011" => y <= "110100000";
					when "11110011100" => y <= "110100001";
					when "11110011101" => y <= "110100010";
					when "11110011110" => y <= "110100011";
					when "11110011111" => y <= "110100100";
					when "11110100000" => y <= "110100101";
					when "11110100001" => y <= "110100110";
					when "11110100010" => y <= "110100111";
					when "11110100011" => y <= "110100111";
					when "11110100100" => y <= "110101000";
					when "11110100101" => y <= "110101001";
					when "11110100110" => y <= "110101010";
					when "11110100111" => y <= "110101011";
					when "11110101000" => y <= "110101100";
					when "11110101001" => y <= "110101101";
					when "11110101010" => y <= "110101110";
					when "11110101011" => y <= "110101110";
					when "11110101100" => y <= "110101111";
					when "11110101101" => y <= "110110000";
					when "11110101110" => y <= "110110001";
					when "11110101111" => y <= "110110010";
					when "11110110000" => y <= "110110011";
					when "11110110001" => y <= "110110100";
					when "11110110010" => y <= "110110101";
					when "11110110011" => y <= "110110110";
					when "11110110100" => y <= "110110111";
					when "11110110101" => y <= "110111000";
					when "11110110110" => y <= "110111000";
					when "11110110111" => y <= "110111001";
					when "11110111000" => y <= "110111010";
					when "11110111001" => y <= "110111011";
					when "11110111010" => y <= "110111100";
					when "11110111011" => y <= "110111101";
					when "11110111100" => y <= "110111110";
					when "11110111101" => y <= "110111111";
					when "11110111110" => y <= "111000000";
					when "11110111111" => y <= "111000001";
					when "11111000000" => y <= "111000010";
					when "11111000001" => y <= "111000011";
					when "11111000010" => y <= "111000100";
					when "11111000011" => y <= "111000101";
					when "11111000100" => y <= "111000110";
					when "11111000101" => y <= "111000111";
					when "11111000110" => y <= "111000111";
					when "11111000111" => y <= "111001000";
					when "11111001000" => y <= "111001001";
					when "11111001001" => y <= "111001010";
					when "11111001010" => y <= "111001011";
					when "11111001011" => y <= "111001100";
					when "11111001100" => y <= "111001101";
					when "11111001101" => y <= "111001110";
					when "11111001110" => y <= "111001111";
					when "11111001111" => y <= "111010000";
					when "11111010000" => y <= "111010001";
					when "11111010001" => y <= "111010010";
					when "11111010010" => y <= "111010011";
					when "11111010011" => y <= "111010100";
					when "11111010100" => y <= "111010101";
					when "11111010101" => y <= "111010110";
					when "11111010110" => y <= "111010111";
					when "11111010111" => y <= "111011000";
					when "11111011000" => y <= "111011001";
					when "11111011001" => y <= "111011010";
					when "11111011010" => y <= "111011011";
					when "11111011011" => y <= "111011100";
					when "11111011100" => y <= "111011101";
					when "11111011101" => y <= "111011110";
					when "11111011110" => y <= "111011111";
					when "11111011111" => y <= "111100000";
					when "11111100000" => y <= "111100001";
					when "11111100001" => y <= "111100010";
					when "11111100010" => y <= "111100011";
					when "11111100011" => y <= "111100100";
					when "11111100100" => y <= "111100101";
					when "11111100101" => y <= "111100110";
					when "11111100110" => y <= "111100111";
					when "11111100111" => y <= "111101000";
					when "11111101000" => y <= "111101001";
					when "11111101001" => y <= "111101010";
					when "11111101010" => y <= "111101011";
					when "11111101011" => y <= "111101100";
					when "11111101100" => y <= "111101101";
					when "11111101101" => y <= "111101110";
					when "11111101110" => y <= "111101111";
					when "11111101111" => y <= "111110000";
					when "11111110000" => y <= "111110001";
					when "11111110001" => y <= "111110010";
					when "11111110010" => y <= "111110011";
					when "11111110011" => y <= "111110100";
					when "11111110100" => y <= "111110101";
					when "11111110101" => y <= "111110110";
					when "11111110110" => y <= "111110111";
					when "11111110111" => y <= "111111000";
					when "11111111000" => y <= "111111001";
					when "11111111001" => y <= "111111010";
					when "11111111010" => y <= "111111011";
					when "11111111011" => y <= "111111100";
					when "11111111100" => y <= "111111101";
					when "11111111101" => y <= "111111110";
					when "11111111110" => y <= "111111111";
					when "11111111111" => y <= "000000000";
					when "00000000000" => y <= "000000000";
					when "00000000001" => y <= "000000000";
					when "00000000010" => y <= "000000001";
					when "00000000011" => y <= "000000010";
					when "00000000100" => y <= "000000011";
					when "00000000101" => y <= "000000100";
					when "00000000110" => y <= "000000101";
					when "00000000111" => y <= "000000110";
					when "00000001000" => y <= "000000111";
					when "00000001001" => y <= "000001000";
					when "00000001010" => y <= "000001001";
					when "00000001011" => y <= "000001010";
					when "00000001100" => y <= "000001011";
					when "00000001101" => y <= "000001100";
					when "00000001110" => y <= "000001101";
					when "00000001111" => y <= "000001110";
					when "00000010000" => y <= "000001111";
					when "00000010001" => y <= "000010000";
					when "00000010010" => y <= "000010001";
					when "00000010011" => y <= "000010010";
					when "00000010100" => y <= "000010011";
					when "00000010101" => y <= "000010100";
					when "00000010110" => y <= "000010101";
					when "00000010111" => y <= "000010110";
					when "00000011000" => y <= "000010111";
					when "00000011001" => y <= "000011000";
					when "00000011010" => y <= "000011001";
					when "00000011011" => y <= "000011010";
					when "00000011100" => y <= "000011011";
					when "00000011101" => y <= "000011100";
					when "00000011110" => y <= "000011101";
					when "00000011111" => y <= "000011110";
					when "00000100000" => y <= "000011111";
					when "00000100001" => y <= "000100000";
					when "00000100010" => y <= "000100001";
					when "00000100011" => y <= "000100010";
					when "00000100100" => y <= "000100011";
					when "00000100101" => y <= "000100100";
					when "00000100110" => y <= "000100101";
					when "00000100111" => y <= "000100110";
					when "00000101000" => y <= "000100111";
					when "00000101001" => y <= "000101000";
					when "00000101010" => y <= "000101001";
					when "00000101011" => y <= "000101010";
					when "00000101100" => y <= "000101011";
					when "00000101101" => y <= "000101100";
					when "00000101110" => y <= "000101101";
					when "00000101111" => y <= "000101110";
					when "00000110000" => y <= "000101111";
					when "00000110001" => y <= "000110000";
					when "00000110010" => y <= "000110001";
					when "00000110011" => y <= "000110010";
					when "00000110100" => y <= "000110011";
					when "00000110101" => y <= "000110100";
					when "00000110110" => y <= "000110101";
					when "00000110111" => y <= "000110110";
					when "00000111000" => y <= "000110111";
					when "00000111001" => y <= "000111000";
					when "00000111010" => y <= "000111001";
					when "00000111011" => y <= "000111001";
					when "00000111100" => y <= "000111010";
					when "00000111101" => y <= "000111011";
					when "00000111110" => y <= "000111100";
					when "00000111111" => y <= "000111101";
					when "00001000000" => y <= "000111110";
					when "00001000001" => y <= "000111111";
					when "00001000010" => y <= "001000000";
					when "00001000011" => y <= "001000001";
					when "00001000100" => y <= "001000010";
					when "00001000101" => y <= "001000011";
					when "00001000110" => y <= "001000100";
					when "00001000111" => y <= "001000101";
					when "00001001000" => y <= "001000110";
					when "00001001001" => y <= "001000111";
					when "00001001010" => y <= "001001000";
					when "00001001011" => y <= "001001000";
					when "00001001100" => y <= "001001001";
					when "00001001101" => y <= "001001010";
					when "00001001110" => y <= "001001011";
					when "00001001111" => y <= "001001100";
					when "00001010000" => y <= "001001101";
					when "00001010001" => y <= "001001110";
					when "00001010010" => y <= "001001111";
					when "00001010011" => y <= "001010000";
					when "00001010100" => y <= "001010001";
					when "00001010101" => y <= "001010010";
					when "00001010110" => y <= "001010010";
					when "00001010111" => y <= "001010011";
					when "00001011000" => y <= "001010100";
					when "00001011001" => y <= "001010101";
					when "00001011010" => y <= "001010110";
					when "00001011011" => y <= "001010111";
					when "00001011100" => y <= "001011000";
					when "00001011101" => y <= "001011001";
					when "00001011110" => y <= "001011001";
					when "00001011111" => y <= "001011010";
					when "00001100000" => y <= "001011011";
					when "00001100001" => y <= "001011100";
					when "00001100010" => y <= "001011101";
					when "00001100011" => y <= "001011110";
					when "00001100100" => y <= "001011111";
					when "00001100101" => y <= "001100000";
					when "00001100110" => y <= "001100000";
					when "00001100111" => y <= "001100001";
					when "00001101000" => y <= "001100010";
					when "00001101001" => y <= "001100011";
					when "00001101010" => y <= "001100100";
					when "00001101011" => y <= "001100101";
					when "00001101100" => y <= "001100110";
					when "00001101101" => y <= "001100110";
					when "00001101110" => y <= "001100111";
					when "00001101111" => y <= "001101000";
					when "00001110000" => y <= "001101001";
					when "00001110001" => y <= "001101010";
					when "00001110010" => y <= "001101011";
					when "00001110011" => y <= "001101011";
					when "00001110100" => y <= "001101100";
					when "00001110101" => y <= "001101101";
					when "00001110110" => y <= "001101110";
					when "00001110111" => y <= "001101111";
					when "00001111000" => y <= "001101111";
					when "00001111001" => y <= "001110000";
					when "00001111010" => y <= "001110001";
					when "00001111011" => y <= "001110010";
					when "00001111100" => y <= "001110011";
					when "00001111101" => y <= "001110011";
					when "00001111110" => y <= "001110100";
					when "00001111111" => y <= "001110101";
					when "00010000000" => y <= "001110110";
					when "00010000001" => y <= "001110111";
					when "00010000010" => y <= "001110111";
					when "00010000011" => y <= "001111000";
					when "00010000100" => y <= "001111001";
					when "00010000101" => y <= "001111010";
					when "00010000110" => y <= "001111010";
					when "00010000111" => y <= "001111011";
					when "00010001000" => y <= "001111100";
					when "00010001001" => y <= "001111101";
					when "00010001010" => y <= "001111110";
					when "00010001011" => y <= "001111110";
					when "00010001100" => y <= "001111111";
					when "00010001101" => y <= "010000000";
					when "00010001110" => y <= "010000001";
					when "00010001111" => y <= "010000001";
					when "00010010000" => y <= "010000010";
					when "00010010001" => y <= "010000011";
					when "00010010010" => y <= "010000011";
					when "00010010011" => y <= "010000100";
					when "00010010100" => y <= "010000101";
					when "00010010101" => y <= "010000110";
					when "00010010110" => y <= "010000110";
					when "00010010111" => y <= "010000111";
					when "00010011000" => y <= "010001000";
					when "00010011001" => y <= "010001001";
					when "00010011010" => y <= "010001001";
					when "00010011011" => y <= "010001010";
					when "00010011100" => y <= "010001011";
					when "00010011101" => y <= "010001011";
					when "00010011110" => y <= "010001100";
					when "00010011111" => y <= "010001101";
					when "00010100000" => y <= "010001101";
					when "00010100001" => y <= "010001110";
					when "00010100010" => y <= "010001111";
					when "00010100011" => y <= "010010000";
					when "00010100100" => y <= "010010000";
					when "00010100101" => y <= "010010001";
					when "00010100110" => y <= "010010010";
					when "00010100111" => y <= "010010010";
					when "00010101000" => y <= "010010011";
					when "00010101001" => y <= "010010100";
					when "00010101010" => y <= "010010100";
					when "00010101011" => y <= "010010101";
					when "00010101100" => y <= "010010110";
					when "00010101101" => y <= "010010110";
					when "00010101110" => y <= "010010111";
					when "00010101111" => y <= "010011000";
					when "00010110000" => y <= "010011000";
					when "00010110001" => y <= "010011001";
					when "00010110010" => y <= "010011001";
					when "00010110011" => y <= "010011010";
					when "00010110100" => y <= "010011011";
					when "00010110101" => y <= "010011011";
					when "00010110110" => y <= "010011100";
					when "00010110111" => y <= "010011101";
					when "00010111000" => y <= "010011101";
					when "00010111001" => y <= "010011110";
					when "00010111010" => y <= "010011110";
					when "00010111011" => y <= "010011111";
					when "00010111100" => y <= "010100000";
					when "00010111101" => y <= "010100000";
					when "00010111110" => y <= "010100001";
					when "00010111111" => y <= "010100010";
					when "00011000000" => y <= "010100010";
					when "00011000001" => y <= "010100011";
					when "00011000010" => y <= "010100011";
					when "00011000011" => y <= "010100100";
					when "00011000100" => y <= "010100100";
					when "00011000101" => y <= "010100101";
					when "00011000110" => y <= "010100110";
					when "00011000111" => y <= "010100110";
					when "00011001000" => y <= "010100111";
					when "00011001001" => y <= "010100111";
					when "00011001010" => y <= "010101000";
					when "00011001011" => y <= "010101000";
					when "00011001100" => y <= "010101001";
					when "00011001101" => y <= "010101010";
					when "00011001110" => y <= "010101010";
					when "00011001111" => y <= "010101011";
					when "00011010000" => y <= "010101011";
					when "00011010001" => y <= "010101100";
					when "00011010010" => y <= "010101100";
					when "00011010011" => y <= "010101101";
					when "00011010100" => y <= "010101101";
					when "00011010101" => y <= "010101110";
					when "00011010110" => y <= "010101111";
					when "00011010111" => y <= "010101111";
					when "00011011000" => y <= "010110000";
					when "00011011001" => y <= "010110000";
					when "00011011010" => y <= "010110001";
					when "00011011011" => y <= "010110001";
					when "00011011100" => y <= "010110010";
					when "00011011101" => y <= "010110010";
					when "00011011110" => y <= "010110011";
					when "00011011111" => y <= "010110011";
					when "00011100000" => y <= "010110100";
					when "00011100001" => y <= "010110100";
					when "00011100010" => y <= "010110101";
					when "00011100011" => y <= "010110101";
					when "00011100100" => y <= "010110110";
					when "00011100101" => y <= "010110110";
					when "00011100110" => y <= "010110111";
					when "00011100111" => y <= "010110111";
					when "00011101000" => y <= "010111000";
					when "00011101001" => y <= "010111000";
					when "00011101010" => y <= "010111001";
					when "00011101011" => y <= "010111001";
					when "00011101100" => y <= "010111010";
					when "00011101101" => y <= "010111010";
					when "00011101110" => y <= "010111010";
					when "00011101111" => y <= "010111011";
					when "00011110000" => y <= "010111011";
					when "00011110001" => y <= "010111100";
					when "00011110010" => y <= "010111100";
					when "00011110011" => y <= "010111101";
					when "00011110100" => y <= "010111101";
					when "00011110101" => y <= "010111110";
					when "00011110110" => y <= "010111110";
					when "00011110111" => y <= "010111111";
					when "00011111000" => y <= "010111111";
					when "00011111001" => y <= "010111111";
					when "00011111010" => y <= "011000000";
					when "00011111011" => y <= "011000000";
					when "00011111100" => y <= "011000001";
					when "00011111101" => y <= "011000001";
					when "00011111110" => y <= "011000010";
					when "00011111111" => y <= "011000010";
					when "00100000000" => y <= "011000010";
					when "00100000001" => y <= "011000011";
					when "00100000010" => y <= "011000011";
					when "00100000011" => y <= "011000100";
					when "00100000100" => y <= "011000100";
					when "00100000101" => y <= "011000101";
					when "00100000110" => y <= "011000101";
					when "00100000111" => y <= "011000101";
					when "00100001000" => y <= "011000110";
					when "00100001001" => y <= "011000110";
					when "00100001010" => y <= "011000111";
					when "00100001011" => y <= "011000111";
					when "00100001100" => y <= "011000111";
					when "00100001101" => y <= "011001000";
					when "00100001110" => y <= "011001000";
					when "00100001111" => y <= "011001000";
					when "00100010000" => y <= "011001001";
					when "00100010001" => y <= "011001001";
					when "00100010010" => y <= "011001010";
					when "00100010011" => y <= "011001010";
					when "00100010100" => y <= "011001010";
					when "00100010101" => y <= "011001011";
					when "00100010110" => y <= "011001011";
					when "00100010111" => y <= "011001011";
					when "00100011000" => y <= "011001100";
					when "00100011001" => y <= "011001100";
					when "00100011010" => y <= "011001101";
					when "00100011011" => y <= "011001101";
					when "00100011100" => y <= "011001101";
					when "00100011101" => y <= "011001110";
					when "00100011110" => y <= "011001110";
					when "00100011111" => y <= "011001110";
					when "00100100000" => y <= "011001111";
					when "00100100001" => y <= "011001111";
					when "00100100010" => y <= "011001111";
					when "00100100011" => y <= "011010000";
					when "00100100100" => y <= "011010000";
					when "00100100101" => y <= "011010000";
					when "00100100110" => y <= "011010001";
					when "00100100111" => y <= "011010001";
					when "00100101000" => y <= "011010001";
					when "00100101001" => y <= "011010010";
					when "00100101010" => y <= "011010010";
					when "00100101011" => y <= "011010010";
					when "00100101100" => y <= "011010011";
					when "00100101101" => y <= "011010011";
					when "00100101110" => y <= "011010011";
					when "00100101111" => y <= "011010100";
					when "00100110000" => y <= "011010100";
					when "00100110001" => y <= "011010100";
					when "00100110010" => y <= "011010101";
					when "00100110011" => y <= "011010101";
					when "00100110100" => y <= "011010101";
					when "00100110101" => y <= "011010101";
					when "00100110110" => y <= "011010110";
					when "00100110111" => y <= "011010110";
					when "00100111000" => y <= "011010110";
					when "00100111001" => y <= "011010111";
					when "00100111010" => y <= "011010111";
					when "00100111011" => y <= "011010111";
					when "00100111100" => y <= "011011000";
					when "00100111101" => y <= "011011000";
					when "00100111110" => y <= "011011000";
					when "00100111111" => y <= "011011000";
					when "00101000000" => y <= "011011001";
					when "00101000001" => y <= "011011001";
					when "00101000010" => y <= "011011001";
					when "00101000011" => y <= "011011001";
					when "00101000100" => y <= "011011010";
					when "00101000101" => y <= "011011010";
					when "00101000110" => y <= "011011010";
					when "00101000111" => y <= "011011011";
					when "00101001000" => y <= "011011011";
					when "00101001001" => y <= "011011011";
					when "00101001010" => y <= "011011011";
					when "00101001011" => y <= "011011100";
					when "00101001100" => y <= "011011100";
					when "00101001101" => y <= "011011100";
					when "00101001110" => y <= "011011100";
					when "00101001111" => y <= "011011101";
					when "00101010000" => y <= "011011101";
					when "00101010001" => y <= "011011101";
					when "00101010010" => y <= "011011101";
					when "00101010011" => y <= "011011110";
					when "00101010100" => y <= "011011110";
					when "00101010101" => y <= "011011110";
					when "00101010110" => y <= "011011110";
					when "00101010111" => y <= "011011111";
					when "00101011000" => y <= "011011111";
					when "00101011001" => y <= "011011111";
					when "00101011010" => y <= "011011111";
					when "00101011011" => y <= "011100000";
					when "00101011100" => y <= "011100000";
					when "00101011101" => y <= "011100000";
					when "00101011110" => y <= "011100000";
					when "00101011111" => y <= "011100001";
					when "00101100000" => y <= "011100001";
					when "00101100001" => y <= "011100001";
					when "00101100010" => y <= "011100001";
					when "00101100011" => y <= "011100001";
					when "00101100100" => y <= "011100010";
					when "00101100101" => y <= "011100010";
					when "00101100110" => y <= "011100010";
					when "00101100111" => y <= "011100010";
					when "00101101000" => y <= "011100010";
					when "00101101001" => y <= "011100011";
					when "00101101010" => y <= "011100011";
					when "00101101011" => y <= "011100011";
					when "00101101100" => y <= "011100011";
					when "00101101101" => y <= "011100100";
					when "00101101110" => y <= "011100100";
					when "00101101111" => y <= "011100100";
					when "00101110000" => y <= "011100100";
					when "00101110001" => y <= "011100100";
					when "00101110010" => y <= "011100101";
					when "00101110011" => y <= "011100101";
					when "00101110100" => y <= "011100101";
					when "00101110101" => y <= "011100101";
					when "00101110110" => y <= "011100101";
					when "00101110111" => y <= "011100110";
					when "00101111000" => y <= "011100110";
					when "00101111001" => y <= "011100110";
					when "00101111010" => y <= "011100110";
					when "00101111011" => y <= "011100110";
					when "00101111100" => y <= "011100110";
					when "00101111101" => y <= "011100111";
					when "00101111110" => y <= "011100111";
					when "00101111111" => y <= "011100111";
					when "00110000000" => y <= "011100111";
					when "00110000001" => y <= "011100111";
					when "00110000010" => y <= "011101000";
					when "00110000011" => y <= "011101000";
					when "00110000100" => y <= "011101000";
					when "00110000101" => y <= "011101000";
					when "00110000110" => y <= "011101000";
					when "00110000111" => y <= "011101000";
					when "00110001000" => y <= "011101001";
					when "00110001001" => y <= "011101001";
					when "00110001010" => y <= "011101001";
					when "00110001011" => y <= "011101001";
					when "00110001100" => y <= "011101001";
					when "00110001101" => y <= "011101001";
					when "00110001110" => y <= "011101010";
					when "00110001111" => y <= "011101010";
					when "00110010000" => y <= "011101010";
					when "00110010001" => y <= "011101010";
					when "00110010010" => y <= "011101010";
					when "00110010011" => y <= "011101010";
					when "00110010100" => y <= "011101011";
					when "00110010101" => y <= "011101011";
					when "00110010110" => y <= "011101011";
					when "00110010111" => y <= "011101011";
					when "00110011000" => y <= "011101011";
					when "00110011001" => y <= "011101011";
					when "00110011010" => y <= "011101100";
					when "00110011011" => y <= "011101100";
					when "00110011100" => y <= "011101100";
					when "00110011101" => y <= "011101100";
					when "00110011110" => y <= "011101100";
					when "00110011111" => y <= "011101100";
					when "00110100000" => y <= "011101100";
					when "00110100001" => y <= "011101101";
					when "00110100010" => y <= "011101101";
					when "00110100011" => y <= "011101101";
					when "00110100100" => y <= "011101101";
					when "00110100101" => y <= "011101101";
					when "00110100110" => y <= "011101101";
					when "00110100111" => y <= "011101101";
					when "00110101000" => y <= "011101110";
					when "00110101001" => y <= "011101110";
					when "00110101010" => y <= "011101110";
					when "00110101011" => y <= "011101110";
					when "00110101100" => y <= "011101110";
					when "00110101101" => y <= "011101110";
					when "00110101110" => y <= "011101110";
					when "00110101111" => y <= "011101110";
					when "00110110000" => y <= "011101111";
					when "00110110001" => y <= "011101111";
					when "00110110010" => y <= "011101111";
					when "00110110011" => y <= "011101111";
					when "00110110100" => y <= "011101111";
					when "00110110101" => y <= "011101111";
					when "00110110110" => y <= "011101111";
					when "00110110111" => y <= "011101111";
					when "00110111000" => y <= "011110000";
					when "00110111001" => y <= "011110000";
					when "00110111010" => y <= "011110000";
					when "00110111011" => y <= "011110000";
					when "00110111100" => y <= "011110000";
					when "00110111101" => y <= "011110000";
					when "00110111110" => y <= "011110000";
					when "00110111111" => y <= "011110000";
					when "00111000000" => y <= "011110000";
					when "00111000001" => y <= "011110001";
					when "00111000010" => y <= "011110001";
					when "00111000011" => y <= "011110001";
					when "00111000100" => y <= "011110001";
					when "00111000101" => y <= "011110001";
					when "00111000110" => y <= "011110001";
					when "00111000111" => y <= "011110001";
					when "00111001000" => y <= "011110001";
					when "00111001001" => y <= "011110001";
					when "00111001010" => y <= "011110010";
					when "00111001011" => y <= "011110010";
					when "00111001100" => y <= "011110010";
					when "00111001101" => y <= "011110010";
					when "00111001110" => y <= "011110010";
					when "00111001111" => y <= "011110010";
					when "00111010000" => y <= "011110010";
					when "00111010001" => y <= "011110010";
					when "00111010010" => y <= "011110010";
					when "00111010011" => y <= "011110011";
					when "00111010100" => y <= "011110011";
					when "00111010101" => y <= "011110011";
					when "00111010110" => y <= "011110011";
					when "00111010111" => y <= "011110011";
					when "00111011000" => y <= "011110011";
					when "00111011001" => y <= "011110011";
					when "00111011010" => y <= "011110011";
					when "00111011011" => y <= "011110011";
					when "00111011100" => y <= "011110011";
					when "00111011101" => y <= "011110011";
					when "00111011110" => y <= "011110100";
					when "00111011111" => y <= "011110100";
					when "00111100000" => y <= "011110100";
					when "00111100001" => y <= "011110100";
					when "00111100010" => y <= "011110100";
					when "00111100011" => y <= "011110100";
					when "00111100100" => y <= "011110100";
					when "00111100101" => y <= "011110100";
					when "00111100110" => y <= "011110100";
					when "00111100111" => y <= "011110100";
					when "00111101000" => y <= "011110100";
					when "00111101001" => y <= "011110101";
					when "00111101010" => y <= "011110101";
					when "00111101011" => y <= "011110101";
					when "00111101100" => y <= "011110101";
					when "00111101101" => y <= "011110101";
					when "00111101110" => y <= "011110101";
					when "00111101111" => y <= "011110101";
					when "00111110000" => y <= "011110101";
					when "00111110001" => y <= "011110101";
					when "00111110010" => y <= "011110101";
					when "00111110011" => y <= "011110101";
					when "00111110100" => y <= "011110101";
					when "00111110101" => y <= "011110101";
					when "00111110110" => y <= "011110110";
					when "00111110111" => y <= "011110110";
					when "00111111000" => y <= "011110110";
					when "00111111001" => y <= "011110110";
					when "00111111010" => y <= "011110110";
					when "00111111011" => y <= "011110110";
					when "00111111100" => y <= "011110110";
					when "00111111101" => y <= "011110110";
					when "00111111110" => y <= "011110110";
					when "00111111111" => y <= "011110110";
					when "01000000000" => y <= "011110110";
					when "01000000001" => y <= "011110110";
					when "01000000010" => y <= "011110110";
					when "01000000011" => y <= "011110111";
					when "01000000100" => y <= "011110111";
					when "01000000101" => y <= "011110111";
					when "01000000110" => y <= "011110111";
					when "01000000111" => y <= "011110111";
					when "01000001000" => y <= "011110111";
					when "01000001001" => y <= "011110111";
					when "01000001010" => y <= "011110111";
					when "01000001011" => y <= "011110111";
					when "01000001100" => y <= "011110111";
					when "01000001101" => y <= "011110111";
					when "01000001110" => y <= "011110111";
					when "01000001111" => y <= "011110111";
					when "01000010000" => y <= "011110111";
					when "01000010001" => y <= "011110111";
					when "01000010010" => y <= "011110111";
					when "01000010011" => y <= "011111000";
					when "01000010100" => y <= "011111000";
					when "01000010101" => y <= "011111000";
					when "01000010110" => y <= "011111000";
					when "01000010111" => y <= "011111000";
					when "01000011000" => y <= "011111000";
					when "01000011001" => y <= "011111000";
					when "01000011010" => y <= "011111000";
					when "01000011011" => y <= "011111000";
					when "01000011100" => y <= "011111000";
					when "01000011101" => y <= "011111000";
					when "01000011110" => y <= "011111000";
					when "01000011111" => y <= "011111000";
					when "01000100000" => y <= "011111000";
					when "01000100001" => y <= "011111000";
					when "01000100010" => y <= "011111000";
					when "01000100011" => y <= "011111000";
					when "01000100100" => y <= "011111001";
					when "01000100101" => y <= "011111001";
					when "01000100110" => y <= "011111001";
					when "01000100111" => y <= "011111001";
					when "01000101000" => y <= "011111001";
					when "01000101001" => y <= "011111001";
					when "01000101010" => y <= "011111001";
					when "01000101011" => y <= "011111001";
					when "01000101100" => y <= "011111001";
					when "01000101101" => y <= "011111001";
					when "01000101110" => y <= "011111001";
					when "01000101111" => y <= "011111001";
					when "01000110000" => y <= "011111001";
					when "01000110001" => y <= "011111001";
					when "01000110010" => y <= "011111001";
					when "01000110011" => y <= "011111001";
					when "01000110100" => y <= "011111001";
					when "01000110101" => y <= "011111001";
					when "01000110110" => y <= "011111001";
					when "01000110111" => y <= "011111001";
					when "01000111000" => y <= "011111010";
					when "01000111001" => y <= "011111010";
					when "01000111010" => y <= "011111010";
					when "01000111011" => y <= "011111010";
					when "01000111100" => y <= "011111010";
					when "01000111101" => y <= "011111010";
					when "01000111110" => y <= "011111010";
					when "01000111111" => y <= "011111010";
					when "01001000000" => y <= "011111010";
					when "01001000001" => y <= "011111010";
					when "01001000010" => y <= "011111010";
					when "01001000011" => y <= "011111010";
					when "01001000100" => y <= "011111010";
					when "01001000101" => y <= "011111010";
					when "01001000110" => y <= "011111010";
					when "01001000111" => y <= "011111010";
					when "01001001000" => y <= "011111010";
					when "01001001001" => y <= "011111010";
					when "01001001010" => y <= "011111010";
					when "01001001011" => y <= "011111010";
					when "01001001100" => y <= "011111010";
					when "01001001101" => y <= "011111010";
					when "01001001110" => y <= "011111010";
					when "01001001111" => y <= "011111010";
					when "01001010000" => y <= "011111011";
					when "01001010001" => y <= "011111011";
					when "01001010010" => y <= "011111011";
					when "01001010011" => y <= "011111011";
					when "01001010100" => y <= "011111011";
					when "01001010101" => y <= "011111011";
					when "01001010110" => y <= "011111011";
					when "01001010111" => y <= "011111011";
					when "01001011000" => y <= "011111011";
					when "01001011001" => y <= "011111011";
					when "01001011010" => y <= "011111011";
					when "01001011011" => y <= "011111011";
					when "01001011100" => y <= "011111011";
					when "01001011101" => y <= "011111011";
					when "01001011110" => y <= "011111011";
					when "01001011111" => y <= "011111011";
					when "01001100000" => y <= "011111011";
					when "01001100001" => y <= "011111011";
					when "01001100010" => y <= "011111011";
					when "01001100011" => y <= "011111011";
					when "01001100100" => y <= "011111011";
					when "01001100101" => y <= "011111011";
					when "01001100110" => y <= "011111011";
					when "01001100111" => y <= "011111011";
					when "01001101000" => y <= "011111011";
					when "01001101001" => y <= "011111011";
					when "01001101010" => y <= "011111011";
					when "01001101011" => y <= "011111011";
					when "01001101100" => y <= "011111011";
					when "01001101101" => y <= "011111100";
					when "01001101110" => y <= "011111100";
					when "01001101111" => y <= "011111100";
					when "01001110000" => y <= "011111100";
					when "01001110001" => y <= "011111100";
					when "01001110010" => y <= "011111100";
					when "01001110011" => y <= "011111100";
					when "01001110100" => y <= "011111100";
					when "01001110101" => y <= "011111100";
					when "01001110110" => y <= "011111100";
					when "01001110111" => y <= "011111100";
					when "01001111000" => y <= "011111100";
					when "01001111001" => y <= "011111100";
					when "01001111010" => y <= "011111100";
					when "01001111011" => y <= "011111100";
					when "01001111100" => y <= "011111100";
					when "01001111101" => y <= "011111100";
					when "01001111110" => y <= "011111100";
					when "01001111111" => y <= "011111100";
					when "01010000000" => y <= "011111100";
					when "01010000001" => y <= "011111100";
					when "01010000010" => y <= "011111100";
					when "01010000011" => y <= "011111100";
					when "01010000100" => y <= "011111100";
					when "01010000101" => y <= "011111100";
					when "01010000110" => y <= "011111100";
					when "01010000111" => y <= "011111100";
					when "01010001000" => y <= "011111100";
					when "01010001001" => y <= "011111100";
					when "01010001010" => y <= "011111100";
					when "01010001011" => y <= "011111100";
					when "01010001100" => y <= "011111100";
					when "01010001101" => y <= "011111100";
					when "01010001110" => y <= "011111100";
					when "01010001111" => y <= "011111100";
					when "01010010000" => y <= "011111100";
					when "01010010001" => y <= "011111100";
					when "01010010010" => y <= "011111101";
					when "01010010011" => y <= "011111101";
					when "01010010100" => y <= "011111101";
					when "01010010101" => y <= "011111101";
					when "01010010110" => y <= "011111101";
					when "01010010111" => y <= "011111101";
					when "01010011000" => y <= "011111101";
					when "01010011001" => y <= "011111101";
					when "01010011010" => y <= "011111101";
					when "01010011011" => y <= "011111101";
					when "01010011100" => y <= "011111101";
					when "01010011101" => y <= "011111101";
					when "01010011110" => y <= "011111101";
					when "01010011111" => y <= "011111101";
					when "01010100000" => y <= "011111101";
					when "01010100001" => y <= "011111101";
					when "01010100010" => y <= "011111101";
					when "01010100011" => y <= "011111101";
					when "01010100100" => y <= "011111101";
					when "01010100101" => y <= "011111101";
					when "01010100110" => y <= "011111101";
					when "01010100111" => y <= "011111101";
					when "01010101000" => y <= "011111101";
					when "01010101001" => y <= "011111101";
					when "01010101010" => y <= "011111101";
					when "01010101011" => y <= "011111101";
					when "01010101100" => y <= "011111101";
					when "01010101101" => y <= "011111101";
					when "01010101110" => y <= "011111101";
					when "01010101111" => y <= "011111101";
					when "01010110000" => y <= "011111101";
					when "01010110001" => y <= "011111101";
					when "01010110010" => y <= "011111101";
					when "01010110011" => y <= "011111101";
					when "01010110100" => y <= "011111101";
					when "01010110101" => y <= "011111101";
					when "01010110110" => y <= "011111101";
					when "01010110111" => y <= "011111101";
					when "01010111000" => y <= "011111101";
					when "01010111001" => y <= "011111101";
					when "01010111010" => y <= "011111101";
					when "01010111011" => y <= "011111101";
					when "01010111100" => y <= "011111101";
					when "01010111101" => y <= "011111101";
					when "01010111110" => y <= "011111101";
					when "01010111111" => y <= "011111101";
					when "01011000000" => y <= "011111101";
					when "01011000001" => y <= "011111101";
					when "01011000010" => y <= "011111101";
					when "01011000011" => y <= "011111101";
					when "01011000100" => y <= "011111101";
					when "01011000101" => y <= "011111101";
					when "01011000110" => y <= "011111110";
					when "01011000111" => y <= "011111110";
					when "01011001000" => y <= "011111110";
					when "01011001001" => y <= "011111110";
					when "01011001010" => y <= "011111110";
					when "01011001011" => y <= "011111110";
					when "01011001100" => y <= "011111110";
					when "01011001101" => y <= "011111110";
					when "01011001110" => y <= "011111110";
					when "01011001111" => y <= "011111110";
					when "01011010000" => y <= "011111110";
					when "01011010001" => y <= "011111110";
					when "01011010010" => y <= "011111110";
					when "01011010011" => y <= "011111110";
					when "01011010100" => y <= "011111110";
					when "01011010101" => y <= "011111110";
					when "01011010110" => y <= "011111110";
					when "01011010111" => y <= "011111110";
					when "01011011000" => y <= "011111110";
					when "01011011001" => y <= "011111110";
					when "01011011010" => y <= "011111110";
					when "01011011011" => y <= "011111110";
					when "01011011100" => y <= "011111110";
					when "01011011101" => y <= "011111110";
					when "01011011110" => y <= "011111110";
					when "01011011111" => y <= "011111110";
					when "01011100000" => y <= "011111110";
					when "01011100001" => y <= "011111110";
					when "01011100010" => y <= "011111110";
					when "01011100011" => y <= "011111110";
					when "01011100100" => y <= "011111110";
					when "01011100101" => y <= "011111110";
					when "01011100110" => y <= "011111110";
					when "01011100111" => y <= "011111110";
					when "01011101000" => y <= "011111110";
					when "01011101001" => y <= "011111110";
					when "01011101010" => y <= "011111110";
					when "01011101011" => y <= "011111110";
					when "01011101100" => y <= "011111110";
					when "01011101101" => y <= "011111110";
					when "01011101110" => y <= "011111110";
					when "01011101111" => y <= "011111110";
					when "01011110000" => y <= "011111110";
					when "01011110001" => y <= "011111110";
					when "01011110010" => y <= "011111110";
					when "01011110011" => y <= "011111110";
					when "01011110100" => y <= "011111110";
					when "01011110101" => y <= "011111110";
					when "01011110110" => y <= "011111110";
					when "01011110111" => y <= "011111110";
					when "01011111000" => y <= "011111110";
					when "01011111001" => y <= "011111110";
					when "01011111010" => y <= "011111110";
					when "01011111011" => y <= "011111110";
					when "01011111100" => y <= "011111110";
					when "01011111101" => y <= "011111110";
					when "01011111110" => y <= "011111110";
					when "01011111111" => y <= "011111110";
					when others => y <= "011111111";
				end case;
			end if;
		end if;
	end process transfer;
	
	eop <= '1' when load = '1' else '0';

end architecture transfer_function_behaviour;